module gamelogic(input logic clk, input logic rst_n, input logic hit
                input logic stand);



endmodule: gamelogic