module lfsr(input logic clk, input logic rst_n, output logic rand);
    
endmodule: lfsr